-- megafunction wizard: %LPM_ADD_SUB%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_ADD_SUB 

-- ============================================================
-- File Name: megaddsub.vhd
-- Megafunction Name(s):
-- 			LPM_ADD_SUB
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2020  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY lpm;
USE lpm.lpm_components.all;
ENTITY megaddsub IS
 PORT ( add_sub : IN STD_LOGIC ;
 dataa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
 datab : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
 result : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
 overflow : OUT STD_LOGIC );
END megaddsub;
ARCHITECTURE SYN OF megaddsub IS
 SIGNAL sub_wire0 : STD_LOGIC ;
 SIGNAL sub_wire1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
 COMPONENT lpm_add_sub
 GENERIC ( lpm_width : NATURAL;
 lpm_direction : STRING;
 lpm_type : STRING;
 lpm_hint : STRING );
 PORT ( dataa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
 add_sub : IN STD_LOGIC ;
 datab : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
 overflow : OUT STD_LOGIC ;
 result : OUT STD_LOGIC_VECTOR (15 DOWNTO 0) );
 END COMPONENT;
BEGIN
 overflow <= sub_wire0;
 result <= sub_wire1(15 DOWNTO 0);
 lpm_add_sub_component : lpm_add_sub
 GENERIC MAP ( lpm_width => 16,
 lpm_direction => "UNUSED",
 lpm_type => "LPM_ADD_SUB",
 lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO" )
 PORT MAP ( dataa => dataa,
 add_sub => add_sub,
 datab => datab,
 overflow => sub_wire0,
 result => sub_wire1 );
END SYN;