LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE cpulib IS

    -- 1. Hardwired Control Unit (ΕΝΗΜΕΡΩΜΕΝΟ)
    COMPONENT hardwired
        PORT (
            ir    : IN  STD_LOGIC_VECTOR(7 DOWNTO 0); -- Πλέον διαβάζει 8 bits
            clock : IN  STD_LOGIC;
            reset : IN  STD_LOGIC;
            z     : IN  STD_LOGIC;
            mOPs  : OUT STD_LOGIC_VECTOR(28 DOWNTO 0) -- 29 bits για BBUS/BLOAD
        );
    END COMPONENT;

    -- 2. Data Bus (ΕΝΗΜΕΡΩΜΕΝΟ με B Register)
    COMPONENT data_bus
        PORT (
            pc_out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            dr_out, tr_out, r_out, ac_out, mem_out : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            b_out : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- ΝΕΟ: Έξοδος B
            
            pcbus, drbus, trbus, rbus, acbus, membus, busmem : IN STD_LOGIC;
            bbus : IN STD_LOGIC; -- ΝΕΟ: Ενεργοποίηση B Bus
            
            dbus        : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            mem_data_in : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
        );
    END COMPONENT;

    -- 3. ALU Controller (Δεν αλλάζει)
    COMPONENT alus
        PORT (
            rbus, acload, zload, andop    : IN  std_logic;
            orop, notop, xorop, aczero    : IN  std_logic;
            acinc, plus, minus, drbus     : IN  std_logic;
            alus                          : OUT std_logic_vector(6 downto 0)
        );
    END COMPONENT;

    -- 4. Τα υπόλοιπα (Ίδια με πριν)
    COMPONENT regnbit
        GENERIC (n : INTEGER := 8); 
        PORT (din : IN std_logic_vector(n-1 downto 0); clk, rst, ld, inc : IN std_logic; dout : OUT std_logic_vector(n-1 downto 0));
    END COMPONENT;

    COMPONENT alu
        GENERIC (n : INTEGER := 8);
        PORT (ac, db : IN std_logic_vector(n-1 downto 0); alus : IN std_logic_vector(7 downto 1); dout : OUT std_logic_vector(n-1 downto 0); z_out : OUT std_logic);
    END COMPONENT;

    COMPONENT RAM
        PORT (address, data : IN STD_LOGIC_VECTOR(7 DOWNTO 0); clock, wren : IN STD_LOGIC; q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT;

END cpulib;